*Mcgarvey, Sabrina A C4C USAF USAFA CW/CS25           * M c g a r v e y ,   S a b r i n a   A   C 4 C   U S A F   U S A F A   C W / C S 2 5   �F �?X�����F �|X